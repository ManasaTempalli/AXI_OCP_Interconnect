`include "gen_definitions.sv"
`include "gen_macros.sv"
`include "interface.sv"
`include "FIFO.sv"
`include "FIFO_control.sv"

`include "axi_wr_front_end.sv"
`include "axi_rd_front_end.sv"
`include "axi_ocp_converter.sv"

`include "ocp_rd_return_front_end.sv"
`include "ocp_axi_converter.sv"

`include "interconnect.sv"

